//Customed AXIS Master Interface
//
//Interface user logic to axis output
//
//Outsider: Standard AXIS-master Interface
//Insider: DIN_DATA, DIN_VALID, DIN_ACCEP, DIN_TLAST
//
//In my opinion, this is pretty a ugly and redundant design
//the user-in to interface-out has one cycle delay, but 
//again, the relative timing is correct
//
//but it has an internal waiting period, so before all this
//stuff begin to transfer, it will wait for 32 cycles
//during that period, the handshake can't be done, so the 
//reflection is the DIN_ACCEP is always set 0;
`timescale 1 ns / 1 ps
	module axis_bram_adapter_v1_0_M00_AXIS #
	(
		parameter integer C_M_AXIS_TDATA_WIDTH	= 32,
        //what the hell does this interface need to wait 
		parameter integer C_M_START_COUNT	= 32
	)
	(
		// Users to add ports here
		input wire [C_M_AXIS_TDATA_WIDTH-1 : 0] DIN_DATA,
        input wire DIN_VALID,
        input wire DIN_TLAST,
        output wire DIN_ACCEP,//interprete this as internal handshake

		// Global ports
		input wire  M_AXIS_ACLK,
		input wire  M_AXIS_ARESETN,
		// Master Stream Ports. TVALID indicates that the master is driving a valid transfer, A transfer takes place when both TVALID and TREADY are asserted. 
		output wire  M_AXIS_TVALID,
		// TDATA is the primary payload that is used to provide the data that is passing across the interface from the master.
		output wire [C_M_AXIS_TDATA_WIDTH-1 : 0] M_AXIS_TDATA,
		// TSTRB is the byte qualifier that indicates whether the content of the associated byte of TDATA is processed as a data byte or a position byte.
		output wire [(C_M_AXIS_TDATA_WIDTH/8)-1 : 0] M_AXIS_TSTRB,
		// TLAST indicates the boundary of a packet.
		output wire  M_AXIS_TLAST,
		// TREADY indicates that the slave can accept a transfer in the current cycle.
		input wire  M_AXIS_TREADY
	);
	                                                                                     
	// function called clogb2 that returns an integer which has the                      
	// value of the ceiling of the log base 2.                                           
	function integer clogb2 (input integer bit_depth);                                   
	  begin                                                                              
	    for(clogb2=0; bit_depth>0; clogb2=clogb2+1)                                      
	      bit_depth = bit_depth >> 1;                                                    
	  end                                                                                
	endfunction                                                                          
	                                                                                     
	// WAIT_COUNT_BITS is the width of the wait counter.                                 
	localparam integer WAIT_COUNT_BITS = clogb2(C_M_START_COUNT-1);                      
	                                                                                     
	// Define the states of state machine                                                
	// The control state machine oversees the writing of input streaming data to the FIFO,
	// and outputs the streaming data from the FIFO                                      
	parameter [1:0] IDLE = 2'b00,        // This is the initial/idle state               
	                                                                                     
	                INIT_COUNTER  = 2'b01, // This state initializes the counter, once   
	                                // the counter reaches C_M_START_COUNT count,        
	                                // the state machine changes state to SEND_STREAM     
                                    //
	                SEND_STREAM   = 2'b10; // In this state the                          
	                                     // stream data is output through M_AXIS_TDATA   
	// State variable                                                                    
	reg [1:0] mst_exec_state;                                                            
	// AXI Stream internal signals
	//wait counter. The master waits for the user defined number of clock cycles before initiating a transfer.
    reg [WAIT_COUNT_BITS-1: 0]  count;
	//streaming data valid
	wire  	axis_tvalid;
	//streaming data valid delayed by one clock cycle
	reg  	axis_tvalid_delay;
	//Last of the streaming data 
	wire  	axis_tlast;
	//Last of the streaming data delayed by one clock cycle
	reg  	axis_tlast_delay;
	//FIFO implementation signals
	reg [C_M_AXIS_TDATA_WIDTH-1 : 0] stream_data_out;
	wire  	tx_en;
	//The master has issued all the streaming data stored in FIFO
	reg  	tx_done;


	// I/O Connections assignments

	assign M_AXIS_TVALID = axis_tvalid_delay;
	assign M_AXIS_TDATA	= stream_data_out;
	assign M_AXIS_TLAST	= axis_tlast_delay;
	assign M_AXIS_TSTRB	= {(C_M_AXIS_TDATA_WIDTH/8){1'b1}};


    //seems like this stupid fsm start increse its state once power on
    //and only reset at lest at seeing tlast
	always @(posedge M_AXIS_ACLK)                                             
	begin                                                                     
	  if (!M_AXIS_ARESETN)                                                    
	    begin                                                                 
	      mst_exec_state <= IDLE;                                             
	      count    <= 0;                                                      
	    end                                                                   
	  else                                                                    
	    case (mst_exec_state)                                                 
	      IDLE:                                                               
	           mst_exec_state  <= INIT_COUNTER;                              
	                                                                         
	      INIT_COUNTER:                                                       
	       if ( count == C_M_START_COUNT - 1 )                               
	          begin                                                           
	            mst_exec_state  <= SEND_STREAM;                               
	          end                                                             
	        else                                                              
	          begin                                                           
	            count <= count + 1;                                           
	            mst_exec_state  <= INIT_COUNTER;                              
	          end                                                             
	                                                                          
	      SEND_STREAM:                                                        
	       if (tx_done)                                                      
	          begin                                                           
	            mst_exec_state <= IDLE;                                       
	          end                                                             
	        else                                                              
	          begin                                                           
	            mst_exec_state <= SEND_STREAM;                                
	          end                                                             
	    endcase                                                               
	end                                                                       


	assign axis_tvalid = ((mst_exec_state == SEND_STREAM) && DIN_VALID);
	assign axis_tlast = DIN_TLAST; 
	assign tx_en = M_AXIS_TREADY && axis_tvalid;   
    assign DIN_ACCEP = tx_en;

	// Delay the axis_tvalid and axis_tlast signal by one clock cycle                              
	// to match the latency of M_AXIS_TDATA                                                        
    // suppose data, tlast arrive at the sample cycle, and valid is compute 
    // in that cycle as well
	always @(posedge M_AXIS_ACLK)                                                                  
	begin                                                                                          
	  if (!M_AXIS_ARESETN)                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= 1'b0;                                                               
	      axis_tlast_delay <= 1'b0;                                                                
	    end                                                                                        
	  else                                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= axis_tvalid;                                                        
	      axis_tlast_delay <= axis_tlast;                                                          
	    end                                                                                        
	end                                                                                            

    always@(posedge M_AXIS_ACLK)
    begin
        if(!M_AXIS_ARESETN)
        begin
            tx_done <= 1'b0;
        end
        else
        begin
            if(DIN_TLAST)
            begin
                tx_done <= 1'b1;
            end
            else
            begin
                tx_done <= 1'b0;
            end
        end
    end

    // Streaming output data is read from FIFO       
    always @( posedge M_AXIS_ACLK )                  
    begin                                            
      if(!M_AXIS_ARESETN)                            
        begin                                        
          stream_data_out <= 0;                      
        end                                          
      else if (tx_en)  
        begin                                        
          stream_data_out <= DIN_DATA;   
        end                                          
      else
      begin
          stream_data_out <= 0;
      end
    end                                              

endmodule
